132.255.208.0/22
167.249.20.0/22
2803:6780::/32
