2803:9610::/32
